module convolve_window_tb;
	reg signed [15:0] window [0:24];
	reg signed [15:0] filter [0:24];
	reg signed [15:0] value;

    	localparam period = 100;
	
	convolve_window cv(window, filter, value);
	
	initial
	begin
		window = { 
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000,
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000,
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000,
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000
		};
		
		filter = { 
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000,
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000,
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000,
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000
		};

        	#period;

		for (integer i=0; i<25; i++)
		begin
			window[i] = 16'b0000100000000000;
          		filter[i] = 16'b0000100000000000;
		end

        	#period;

		for (integer i=0; i<25; i++)
		begin
				window[i] = 16'b1011000000000000;
          			filter[i] = 16'b0000100000000000;
		end

        	#period;

	end

endmodule
