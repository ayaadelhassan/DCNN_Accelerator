module fortesting(input x,y);





endmodule
