module pool_image_tb;
	reg signed [15:0] image [0:15];
	reg signed [15:0] pooled_image [0:3];

    	localparam period = 100;
	
	pool_image #(.n(4)) pool(image, pooled_image);
	
	initial
	begin
//		image = { 16'b0000010000000000, 16'b0000010000000000, 16'b0000100000000000, 16'b0000110000000000, 
//			16'b0000010000000000, 16'b0000010000000000, 16'b1111110000000000, 16'b1111000000000000,
//			16'b0101000000000000, 16'b0101100000000000, 16'b1011000000000000, 16'b1010100000000000, 
//			16'b0110000000000000, 16'b0110100000000000, 16'b1010000000000000, 16'b1001100000000000
//		};
//		#period;

		image = { 16'b0100010000000000, 16'b0000010100000000, 16'b0100100000000000, 16'b0010110000000000, 
			16'b1100010000000000, 16'b0000010000000000, 16'b1111110011000000, 16'b1111000000000000,
			16'b0101000000000000, 16'b0101100000000000, 16'b1011000000000000, 16'b1010100010000000, 
			16'b0000000000000000, 16'b0110100000000011, 16'b1011000000000000, 16'b1001110000000000
		};
		#period;


	end

endmodule