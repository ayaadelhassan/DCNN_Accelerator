module convolve_image_clked_tb;
	reg signed [15:0] image [0:99];
	reg signed [15:0] filter [0:24];
	reg signed [15:0] convolved_image [0:35];

    	localparam period = 100;
	
	convolve_image #(.n(10)) cv(image, filter, convolved_image);
	
	initial
	begin

        forever begin
        clk = 0;
        #10 clk = ~clk;
        end 
		image = { 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000,
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000,
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000,
			16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000, 16'b0000010000000000
		};
		
		filter = { 
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000,
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000,
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000,
			16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000, 16'b0000100000000000
		};

       	#period;

		for (integer i=0; i<100; i++)
		begin
          		image[i] = 16'b0000010000000000;
		end


		for (integer i=0; i<25; i++)
		begin
          		filter[i] = 16'b0000100000000000;
		end
		
		image[3] = 16'b1010000000000000;
        	
		#period;


	end

endmodule
