/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May  5 19:19:17 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1466647365 */

module Comparitor(Arr0, Arr1, Arr2, Arr3, Arr4, Arr5, Arr6, Arr7, Arr8, Arr9, 
      clk, done, result, enable, reset);
   input [15:0]Arr0;
   input [15:0]Arr1;
   input [15:0]Arr2;
   input [15:0]Arr3;
   input [15:0]Arr4;
   input [15:0]Arr5;
   input [15:0]Arr6;
   input [15:0]Arr7;
   input [15:0]Arr8;
   input [15:0]Arr9;
   input clk;
   output done;
   output [3:0]result;
   input enable;
   input reset;

   wire n_0_0;
   wire n_0_27;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire [15:0]max;
   wire n_0_30;
   wire [3:0]i;
   wire n_0_5;
   wire n_0_0_2;
   wire n_0_0_0;
   wire n_0_0_3;
   wire n_0_0_1;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_0_4;
   wire n_0_31;
   wire n_0_29;
   wire [3:0]maxIndex;
   wire n_0_28;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_32;
   wire n_0_0_33;
   wire n_0_0_34;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_0_41;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_10;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_11;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_12;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_13;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_14;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_15;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_16;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_17;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_18;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_19;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_20;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_21;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_22;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_23;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_24;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_25;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_6;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_26;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;

   CLKGATETST_X1 clk_gate_result_reg (.CK(clk), .E(n_0_26), .SE(1'b0), .GCK(
      n_0_0));
   DFF_X1 \result_reg[3]  (.D(n_0_1), .CK(n_0_0), .Q(result[3]), .QN());
   DFF_X1 \result_reg[2]  (.D(n_0_2), .CK(n_0_0), .Q(result[2]), .QN());
   DFF_X1 \result_reg[1]  (.D(n_0_3), .CK(n_0_0), .Q(result[1]), .QN());
   DFF_X1 \result_reg[0]  (.D(n_0_4), .CK(n_0_0), .Q(result[0]), .QN());
   DFF_X1 done_reg (.D(n_0_27), .CK(clk), .Q(done), .QN());
   MUX2_X1 done_reg_enable_mux_0 (.A(done), .B(n_0_26), .S(n_0_29), .Z(n_0_27));
   DFF_X1 \maxIndex_reg[3]  (.D(maxIndex[3]), .CK(n_0_5), .Q(n_0_1), .QN());
   DFF_X1 \maxIndex_reg[2]  (.D(maxIndex[2]), .CK(n_0_5), .Q(n_0_2), .QN());
   DFF_X1 \maxIndex_reg[1]  (.D(maxIndex[1]), .CK(n_0_5), .Q(n_0_3), .QN());
   DFF_X1 \maxIndex_reg[0]  (.D(maxIndex[0]), .CK(n_0_5), .Q(n_0_4), .QN());
   DFF_X1 \max_reg[15]  (.D(n_0_25), .CK(n_0_5), .Q(max[15]), .QN());
   DFF_X1 \max_reg[14]  (.D(n_0_24), .CK(n_0_5), .Q(max[14]), .QN());
   DFF_X1 \max_reg[13]  (.D(n_0_23), .CK(n_0_5), .Q(max[13]), .QN());
   DFF_X1 \max_reg[12]  (.D(n_0_22), .CK(n_0_5), .Q(max[12]), .QN());
   DFF_X1 \max_reg[11]  (.D(n_0_21), .CK(n_0_5), .Q(max[11]), .QN());
   DFF_X1 \max_reg[10]  (.D(n_0_20), .CK(n_0_5), .Q(max[10]), .QN());
   DFF_X1 \max_reg[9]  (.D(n_0_19), .CK(n_0_5), .Q(max[9]), .QN());
   DFF_X1 \max_reg[8]  (.D(n_0_18), .CK(n_0_5), .Q(max[8]), .QN());
   DFF_X1 \max_reg[7]  (.D(n_0_17), .CK(n_0_5), .Q(max[7]), .QN());
   DFF_X1 \max_reg[6]  (.D(n_0_16), .CK(n_0_5), .Q(max[6]), .QN());
   DFF_X1 \max_reg[5]  (.D(n_0_15), .CK(n_0_5), .Q(max[5]), .QN());
   DFF_X1 \max_reg[4]  (.D(n_0_14), .CK(n_0_5), .Q(max[4]), .QN());
   DFF_X1 \max_reg[3]  (.D(n_0_13), .CK(n_0_5), .Q(max[3]), .QN());
   DFF_X1 \max_reg[2]  (.D(n_0_12), .CK(n_0_5), .Q(max[2]), .QN());
   DFF_X1 \max_reg[1]  (.D(n_0_11), .CK(n_0_5), .Q(max[1]), .QN());
   DFF_X1 \max_reg[0]  (.D(n_0_10), .CK(n_0_5), .Q(max[0]), .QN());
   CLKGATETST_X1 clk_gate_i_reg (.CK(clk), .E(n_0_31), .SE(1'b0), .GCK(n_0_30));
   DFF_X1 \i_reg[3]  (.D(n_0_9), .CK(n_0_30), .Q(i[3]), .QN());
   DFF_X1 \i_reg[2]  (.D(n_0_8), .CK(n_0_30), .Q(i[2]), .QN());
   DFF_X1 \i_reg[1]  (.D(n_0_7), .CK(n_0_30), .Q(i[1]), .QN());
   DFF_X1 \i_reg[0]  (.D(n_0_6), .CK(n_0_30), .Q(i[0]), .QN());
   CLKGATETST_X1 clk_gate_maxIndex_reg (.CK(clk), .E(n_0_28), .SE(1'b0), 
      .GCK(n_0_5));
   HA_X1 i_0_0_0 (.A(i[1]), .B(i[0]), .CO(n_0_0_0), .S(n_0_0_2));
   HA_X1 i_0_0_1 (.A(i[2]), .B(n_0_0_0), .CO(n_0_0_1), .S(n_0_0_3));
   AND2_X1 i_0_0_2 (.A1(n_0_0_2), .A2(n_0_0_323), .ZN(n_0_7));
   AND2_X1 i_0_0_3 (.A1(n_0_0_3), .A2(n_0_0_323), .ZN(n_0_8));
   AOI21_X1 i_0_0_4 (.A(n_0_0_4), .B1(n_0_0_1), .B2(i[3]), .ZN(n_0_9));
   OAI21_X1 i_0_0_5 (.A(n_0_0_323), .B1(n_0_0_1), .B2(i[3]), .ZN(n_0_0_4));
   OR2_X1 i_0_0_6 (.A1(reset), .A2(n_0_0_323), .ZN(n_0_31));
   OR2_X1 i_0_0_7 (.A1(reset), .A2(n_0_26), .ZN(n_0_29));
   AOI21_X1 i_0_0_8 (.A(n_0_6), .B1(n_0_0_325), .B2(i[3]), .ZN(maxIndex[0]));
   NAND3_X1 i_0_0_9 (.A1(n_0_0_130), .A2(n_0_0_54), .A3(n_0_0_5), .ZN(n_0_28));
   AOI22_X1 i_0_0_10 (.A1(n_0_0_314), .A2(n_0_0_30), .B1(n_0_0_6), .B2(n_0_0_316), 
      .ZN(n_0_0_5));
   OAI22_X1 i_0_0_11 (.A1(n_0_0_8), .A2(n_0_0_7), .B1(n_0_0_357), .B2(Arr3[15]), 
      .ZN(n_0_0_6));
   OAI22_X1 i_0_0_12 (.A1(n_0_0_356), .A2(Arr3[14]), .B1(n_0_0_332), .B2(max[15]), 
      .ZN(n_0_0_7));
   AOI21_X1 i_0_0_13 (.A(n_0_0_9), .B1(Arr3[14]), .B2(n_0_0_356), .ZN(n_0_0_8));
   AOI21_X1 i_0_0_14 (.A(n_0_0_29), .B1(n_0_0_11), .B2(n_0_0_10), .ZN(n_0_0_9));
   AOI22_X1 i_0_0_15 (.A1(n_0_0_355), .A2(Arr3[13]), .B1(n_0_0_354), .B2(
      Arr3[12]), .ZN(n_0_0_10));
   OAI221_X1 i_0_0_16 (.A(n_0_0_12), .B1(Arr3[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr3[12]), .ZN(n_0_0_11));
   NAND2_X1 i_0_0_17 (.A1(n_0_0_14), .A2(n_0_0_13), .ZN(n_0_0_12));
   AOI22_X1 i_0_0_18 (.A1(n_0_0_353), .A2(Arr3[11]), .B1(n_0_0_352), .B2(
      Arr3[10]), .ZN(n_0_0_13));
   OAI221_X1 i_0_0_19 (.A(n_0_0_15), .B1(Arr3[9]), .B2(n_0_0_351), .C1(n_0_0_352), 
      .C2(Arr3[10]), .ZN(n_0_0_14));
   NAND2_X1 i_0_0_20 (.A1(n_0_0_17), .A2(n_0_0_16), .ZN(n_0_0_15));
   AOI22_X1 i_0_0_21 (.A1(n_0_0_351), .A2(Arr3[9]), .B1(n_0_0_350), .B2(Arr3[8]), 
      .ZN(n_0_0_16));
   OAI221_X1 i_0_0_22 (.A(n_0_0_18), .B1(Arr3[7]), .B2(n_0_0_349), .C1(n_0_0_350), 
      .C2(Arr3[8]), .ZN(n_0_0_17));
   NAND2_X1 i_0_0_23 (.A1(n_0_0_20), .A2(n_0_0_19), .ZN(n_0_0_18));
   AOI22_X1 i_0_0_24 (.A1(n_0_0_349), .A2(Arr3[7]), .B1(n_0_0_348), .B2(Arr3[6]), 
      .ZN(n_0_0_19));
   OAI221_X1 i_0_0_25 (.A(n_0_0_21), .B1(Arr3[5]), .B2(n_0_0_347), .C1(n_0_0_348), 
      .C2(Arr3[6]), .ZN(n_0_0_20));
   NAND2_X1 i_0_0_26 (.A1(n_0_0_23), .A2(n_0_0_22), .ZN(n_0_0_21));
   AOI22_X1 i_0_0_27 (.A1(n_0_0_347), .A2(Arr3[5]), .B1(n_0_0_346), .B2(Arr3[4]), 
      .ZN(n_0_0_22));
   OAI21_X1 i_0_0_28 (.A(n_0_0_24), .B1(Arr3[4]), .B2(n_0_0_346), .ZN(n_0_0_23));
   OAI21_X1 i_0_0_29 (.A(n_0_0_25), .B1(n_0_0_331), .B2(max[3]), .ZN(n_0_0_24));
   OAI221_X1 i_0_0_30 (.A(n_0_0_26), .B1(Arr3[2]), .B2(n_0_0_344), .C1(n_0_0_345), 
      .C2(Arr3[3]), .ZN(n_0_0_25));
   NAND2_X1 i_0_0_31 (.A1(n_0_0_27), .A2(n_0_0_28), .ZN(n_0_0_26));
   AOI22_X1 i_0_0_32 (.A1(n_0_0_344), .A2(Arr3[2]), .B1(n_0_0_343), .B2(Arr3[1]), 
      .ZN(n_0_0_27));
   OAI211_X1 i_0_0_33 (.A(n_0_0_342), .B(Arr3[0]), .C1(n_0_0_343), .C2(Arr3[1]), 
      .ZN(n_0_0_28));
   NOR2_X1 i_0_0_34 (.A1(n_0_0_355), .A2(Arr3[13]), .ZN(n_0_0_29));
   OAI22_X1 i_0_0_35 (.A1(n_0_0_32), .A2(n_0_0_31), .B1(n_0_0_357), .B2(Arr4[15]), 
      .ZN(n_0_0_30));
   OAI22_X1 i_0_0_36 (.A1(n_0_0_356), .A2(Arr4[14]), .B1(n_0_0_334), .B2(max[15]), 
      .ZN(n_0_0_31));
   AOI21_X1 i_0_0_37 (.A(n_0_0_33), .B1(Arr4[14]), .B2(n_0_0_356), .ZN(n_0_0_32));
   AOI21_X1 i_0_0_38 (.A(n_0_0_53), .B1(n_0_0_35), .B2(n_0_0_34), .ZN(n_0_0_33));
   AOI22_X1 i_0_0_39 (.A1(n_0_0_355), .A2(Arr4[13]), .B1(n_0_0_354), .B2(
      Arr4[12]), .ZN(n_0_0_34));
   OAI221_X1 i_0_0_40 (.A(n_0_0_36), .B1(Arr4[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr4[12]), .ZN(n_0_0_35));
   NAND2_X1 i_0_0_41 (.A1(n_0_0_38), .A2(n_0_0_37), .ZN(n_0_0_36));
   AOI22_X1 i_0_0_42 (.A1(n_0_0_353), .A2(Arr4[11]), .B1(n_0_0_352), .B2(
      Arr4[10]), .ZN(n_0_0_37));
   OAI221_X1 i_0_0_43 (.A(n_0_0_39), .B1(Arr4[9]), .B2(n_0_0_351), .C1(n_0_0_352), 
      .C2(Arr4[10]), .ZN(n_0_0_38));
   NAND2_X1 i_0_0_44 (.A1(n_0_0_41), .A2(n_0_0_40), .ZN(n_0_0_39));
   AOI22_X1 i_0_0_45 (.A1(n_0_0_351), .A2(Arr4[9]), .B1(n_0_0_350), .B2(Arr4[8]), 
      .ZN(n_0_0_40));
   OAI221_X1 i_0_0_46 (.A(n_0_0_42), .B1(Arr4[7]), .B2(n_0_0_349), .C1(n_0_0_350), 
      .C2(Arr4[8]), .ZN(n_0_0_41));
   NAND2_X1 i_0_0_47 (.A1(n_0_0_44), .A2(n_0_0_43), .ZN(n_0_0_42));
   AOI22_X1 i_0_0_48 (.A1(n_0_0_349), .A2(Arr4[7]), .B1(n_0_0_348), .B2(Arr4[6]), 
      .ZN(n_0_0_43));
   OAI221_X1 i_0_0_49 (.A(n_0_0_45), .B1(Arr4[5]), .B2(n_0_0_347), .C1(n_0_0_348), 
      .C2(Arr4[6]), .ZN(n_0_0_44));
   NAND2_X1 i_0_0_50 (.A1(n_0_0_47), .A2(n_0_0_46), .ZN(n_0_0_45));
   AOI22_X1 i_0_0_51 (.A1(n_0_0_347), .A2(Arr4[5]), .B1(n_0_0_346), .B2(Arr4[4]), 
      .ZN(n_0_0_46));
   OAI21_X1 i_0_0_52 (.A(n_0_0_48), .B1(Arr4[4]), .B2(n_0_0_346), .ZN(n_0_0_47));
   OAI21_X1 i_0_0_53 (.A(n_0_0_49), .B1(n_0_0_333), .B2(max[3]), .ZN(n_0_0_48));
   OAI221_X1 i_0_0_54 (.A(n_0_0_50), .B1(Arr4[2]), .B2(n_0_0_344), .C1(n_0_0_345), 
      .C2(Arr4[3]), .ZN(n_0_0_49));
   NAND2_X1 i_0_0_55 (.A1(n_0_0_51), .A2(n_0_0_52), .ZN(n_0_0_50));
   AOI22_X1 i_0_0_56 (.A1(n_0_0_344), .A2(Arr4[2]), .B1(n_0_0_343), .B2(Arr4[1]), 
      .ZN(n_0_0_51));
   OAI211_X1 i_0_0_57 (.A(n_0_0_342), .B(Arr4[0]), .C1(n_0_0_343), .C2(Arr4[1]), 
      .ZN(n_0_0_52));
   NOR2_X1 i_0_0_58 (.A1(n_0_0_355), .A2(Arr4[13]), .ZN(n_0_0_53));
   AND3_X1 i_0_0_59 (.A1(n_0_0_105), .A2(n_0_0_80), .A3(n_0_0_55), .ZN(n_0_0_54));
   NAND3_X1 i_0_0_60 (.A1(n_0_0_57), .A2(n_0_0_56), .A3(n_0_0_309), .ZN(n_0_0_55));
   NAND2_X1 i_0_0_61 (.A1(n_0_0_357), .A2(Arr6[15]), .ZN(n_0_0_56));
   OAI211_X1 i_0_0_62 (.A(n_0_0_59), .B(n_0_0_58), .C1(n_0_0_357), .C2(Arr6[15]), 
      .ZN(n_0_0_57));
   NAND2_X1 i_0_0_63 (.A1(n_0_0_356), .A2(Arr6[14]), .ZN(n_0_0_58));
   OAI221_X1 i_0_0_64 (.A(n_0_0_60), .B1(Arr6[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr6[14]), .ZN(n_0_0_59));
   NAND2_X1 i_0_0_65 (.A1(n_0_0_62), .A2(n_0_0_61), .ZN(n_0_0_60));
   AOI22_X1 i_0_0_66 (.A1(n_0_0_355), .A2(Arr6[13]), .B1(n_0_0_354), .B2(
      Arr6[12]), .ZN(n_0_0_61));
   OAI221_X1 i_0_0_67 (.A(n_0_0_63), .B1(Arr6[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr6[12]), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_68 (.A1(n_0_0_65), .A2(n_0_0_64), .ZN(n_0_0_63));
   AOI22_X1 i_0_0_69 (.A1(n_0_0_353), .A2(Arr6[11]), .B1(n_0_0_352), .B2(
      Arr6[10]), .ZN(n_0_0_64));
   OAI221_X1 i_0_0_70 (.A(n_0_0_66), .B1(Arr6[9]), .B2(n_0_0_351), .C1(n_0_0_352), 
      .C2(Arr6[10]), .ZN(n_0_0_65));
   NAND2_X1 i_0_0_71 (.A1(n_0_0_68), .A2(n_0_0_67), .ZN(n_0_0_66));
   AOI22_X1 i_0_0_72 (.A1(n_0_0_351), .A2(Arr6[9]), .B1(n_0_0_350), .B2(Arr6[8]), 
      .ZN(n_0_0_67));
   OAI221_X1 i_0_0_73 (.A(n_0_0_69), .B1(Arr6[7]), .B2(n_0_0_349), .C1(n_0_0_350), 
      .C2(Arr6[8]), .ZN(n_0_0_68));
   NAND2_X1 i_0_0_74 (.A1(n_0_0_71), .A2(n_0_0_70), .ZN(n_0_0_69));
   AOI22_X1 i_0_0_75 (.A1(n_0_0_349), .A2(Arr6[7]), .B1(n_0_0_348), .B2(Arr6[6]), 
      .ZN(n_0_0_70));
   OAI221_X1 i_0_0_76 (.A(n_0_0_72), .B1(Arr6[5]), .B2(n_0_0_347), .C1(n_0_0_348), 
      .C2(Arr6[6]), .ZN(n_0_0_71));
   NAND2_X1 i_0_0_77 (.A1(n_0_0_74), .A2(n_0_0_73), .ZN(n_0_0_72));
   AOI22_X1 i_0_0_78 (.A1(n_0_0_347), .A2(Arr6[5]), .B1(n_0_0_346), .B2(Arr6[4]), 
      .ZN(n_0_0_73));
   OAI21_X1 i_0_0_79 (.A(n_0_0_75), .B1(Arr6[4]), .B2(n_0_0_346), .ZN(n_0_0_74));
   OAI21_X1 i_0_0_80 (.A(n_0_0_76), .B1(n_0_0_337), .B2(max[3]), .ZN(n_0_0_75));
   OAI221_X1 i_0_0_81 (.A(n_0_0_77), .B1(Arr6[2]), .B2(n_0_0_344), .C1(n_0_0_345), 
      .C2(Arr6[3]), .ZN(n_0_0_76));
   NAND2_X1 i_0_0_82 (.A1(n_0_0_78), .A2(n_0_0_79), .ZN(n_0_0_77));
   AOI22_X1 i_0_0_83 (.A1(n_0_0_344), .A2(Arr6[2]), .B1(n_0_0_343), .B2(Arr6[1]), 
      .ZN(n_0_0_78));
   OAI211_X1 i_0_0_84 (.A(n_0_0_342), .B(Arr6[0]), .C1(n_0_0_343), .C2(Arr6[1]), 
      .ZN(n_0_0_79));
   NAND3_X1 i_0_0_85 (.A1(n_0_0_82), .A2(n_0_0_81), .A3(n_0_0_307), .ZN(n_0_0_80));
   NAND2_X1 i_0_0_86 (.A1(n_0_0_357), .A2(Arr1[15]), .ZN(n_0_0_81));
   OAI211_X1 i_0_0_87 (.A(n_0_0_84), .B(n_0_0_83), .C1(n_0_0_357), .C2(Arr1[15]), 
      .ZN(n_0_0_82));
   NAND2_X1 i_0_0_88 (.A1(n_0_0_356), .A2(Arr1[14]), .ZN(n_0_0_83));
   OAI221_X1 i_0_0_89 (.A(n_0_0_85), .B1(Arr1[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr1[14]), .ZN(n_0_0_84));
   NAND2_X1 i_0_0_90 (.A1(n_0_0_87), .A2(n_0_0_86), .ZN(n_0_0_85));
   AOI22_X1 i_0_0_91 (.A1(n_0_0_355), .A2(Arr1[13]), .B1(n_0_0_354), .B2(
      Arr1[12]), .ZN(n_0_0_86));
   OAI221_X1 i_0_0_92 (.A(n_0_0_88), .B1(Arr1[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr1[12]), .ZN(n_0_0_87));
   NAND2_X1 i_0_0_93 (.A1(n_0_0_90), .A2(n_0_0_89), .ZN(n_0_0_88));
   AOI22_X1 i_0_0_94 (.A1(n_0_0_353), .A2(Arr1[11]), .B1(n_0_0_352), .B2(
      Arr1[10]), .ZN(n_0_0_89));
   OAI21_X1 i_0_0_95 (.A(n_0_0_91), .B1(Arr1[10]), .B2(n_0_0_352), .ZN(n_0_0_90));
   OAI21_X1 i_0_0_96 (.A(n_0_0_92), .B1(n_0_0_328), .B2(max[9]), .ZN(n_0_0_91));
   OAI221_X1 i_0_0_97 (.A(n_0_0_93), .B1(Arr1[8]), .B2(n_0_0_350), .C1(n_0_0_351), 
      .C2(Arr1[9]), .ZN(n_0_0_92));
   NAND2_X1 i_0_0_98 (.A1(n_0_0_95), .A2(n_0_0_94), .ZN(n_0_0_93));
   AOI22_X1 i_0_0_99 (.A1(n_0_0_350), .A2(Arr1[8]), .B1(n_0_0_349), .B2(Arr1[7]), 
      .ZN(n_0_0_94));
   OAI221_X1 i_0_0_100 (.A(n_0_0_96), .B1(Arr1[6]), .B2(n_0_0_348), .C1(
      n_0_0_349), .C2(Arr1[7]), .ZN(n_0_0_95));
   NAND2_X1 i_0_0_101 (.A1(n_0_0_98), .A2(n_0_0_97), .ZN(n_0_0_96));
   AOI22_X1 i_0_0_102 (.A1(n_0_0_348), .A2(Arr1[6]), .B1(n_0_0_347), .B2(Arr1[5]), 
      .ZN(n_0_0_97));
   OAI221_X1 i_0_0_103 (.A(n_0_0_99), .B1(Arr1[4]), .B2(n_0_0_346), .C1(
      n_0_0_347), .C2(Arr1[5]), .ZN(n_0_0_98));
   NAND2_X1 i_0_0_104 (.A1(n_0_0_101), .A2(n_0_0_100), .ZN(n_0_0_99));
   AOI22_X1 i_0_0_105 (.A1(n_0_0_346), .A2(Arr1[4]), .B1(n_0_0_345), .B2(Arr1[3]), 
      .ZN(n_0_0_100));
   OAI221_X1 i_0_0_106 (.A(n_0_0_102), .B1(Arr1[2]), .B2(n_0_0_344), .C1(
      n_0_0_345), .C2(Arr1[3]), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_107 (.A1(n_0_0_103), .A2(n_0_0_104), .ZN(n_0_0_102));
   AOI22_X1 i_0_0_108 (.A1(n_0_0_344), .A2(Arr1[2]), .B1(n_0_0_343), .B2(Arr1[1]), 
      .ZN(n_0_0_103));
   OAI211_X1 i_0_0_109 (.A(n_0_0_342), .B(Arr1[0]), .C1(n_0_0_343), .C2(Arr1[1]), 
      .ZN(n_0_0_104));
   AOI21_X1 i_0_0_110 (.A(n_0_0_106), .B1(n_0_0_313), .B2(reset), .ZN(n_0_0_105));
   AOI21_X1 i_0_0_111 (.A(n_0_0_107), .B1(n_0_0_109), .B2(n_0_0_108), .ZN(
      n_0_0_106));
   OAI21_X1 i_0_0_112 (.A(n_0_0_310), .B1(n_0_0_336), .B2(max[15]), .ZN(
      n_0_0_107));
   AOI22_X1 i_0_0_113 (.A1(n_0_0_356), .A2(Arr5[14]), .B1(n_0_0_336), .B2(
      max[15]), .ZN(n_0_0_108));
   OAI221_X1 i_0_0_114 (.A(n_0_0_110), .B1(Arr5[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr5[14]), .ZN(n_0_0_109));
   NAND2_X1 i_0_0_115 (.A1(n_0_0_112), .A2(n_0_0_111), .ZN(n_0_0_110));
   AOI22_X1 i_0_0_116 (.A1(n_0_0_355), .A2(Arr5[13]), .B1(n_0_0_354), .B2(
      Arr5[12]), .ZN(n_0_0_111));
   OAI221_X1 i_0_0_117 (.A(n_0_0_113), .B1(Arr5[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr5[12]), .ZN(n_0_0_112));
   NAND2_X1 i_0_0_118 (.A1(n_0_0_115), .A2(n_0_0_114), .ZN(n_0_0_113));
   AOI22_X1 i_0_0_119 (.A1(n_0_0_353), .A2(Arr5[11]), .B1(n_0_0_352), .B2(
      Arr5[10]), .ZN(n_0_0_114));
   OAI221_X1 i_0_0_120 (.A(n_0_0_116), .B1(Arr5[9]), .B2(n_0_0_351), .C1(
      n_0_0_352), .C2(Arr5[10]), .ZN(n_0_0_115));
   NAND2_X1 i_0_0_121 (.A1(n_0_0_118), .A2(n_0_0_117), .ZN(n_0_0_116));
   AOI22_X1 i_0_0_122 (.A1(n_0_0_351), .A2(Arr5[9]), .B1(n_0_0_350), .B2(Arr5[8]), 
      .ZN(n_0_0_117));
   OAI21_X1 i_0_0_123 (.A(n_0_0_119), .B1(Arr5[8]), .B2(n_0_0_350), .ZN(
      n_0_0_118));
   OAI21_X1 i_0_0_124 (.A(n_0_0_120), .B1(n_0_0_335), .B2(max[7]), .ZN(n_0_0_119));
   OAI221_X1 i_0_0_125 (.A(n_0_0_121), .B1(Arr5[6]), .B2(n_0_0_348), .C1(
      n_0_0_349), .C2(Arr5[7]), .ZN(n_0_0_120));
   NAND2_X1 i_0_0_126 (.A1(n_0_0_123), .A2(n_0_0_122), .ZN(n_0_0_121));
   AOI22_X1 i_0_0_127 (.A1(n_0_0_348), .A2(Arr5[6]), .B1(n_0_0_347), .B2(Arr5[5]), 
      .ZN(n_0_0_122));
   OAI221_X1 i_0_0_128 (.A(n_0_0_124), .B1(Arr5[4]), .B2(n_0_0_346), .C1(
      n_0_0_347), .C2(Arr5[5]), .ZN(n_0_0_123));
   NAND2_X1 i_0_0_129 (.A1(n_0_0_126), .A2(n_0_0_125), .ZN(n_0_0_124));
   AOI22_X1 i_0_0_130 (.A1(n_0_0_346), .A2(Arr5[4]), .B1(n_0_0_345), .B2(Arr5[3]), 
      .ZN(n_0_0_125));
   OAI221_X1 i_0_0_131 (.A(n_0_0_127), .B1(Arr5[2]), .B2(n_0_0_344), .C1(
      n_0_0_345), .C2(Arr5[3]), .ZN(n_0_0_126));
   NAND2_X1 i_0_0_132 (.A1(n_0_0_128), .A2(n_0_0_129), .ZN(n_0_0_127));
   AOI22_X1 i_0_0_133 (.A1(n_0_0_344), .A2(Arr5[2]), .B1(n_0_0_343), .B2(Arr5[1]), 
      .ZN(n_0_0_128));
   OAI211_X1 i_0_0_134 (.A(n_0_0_342), .B(Arr5[0]), .C1(n_0_0_343), .C2(Arr5[1]), 
      .ZN(n_0_0_129));
   NOR4_X1 i_0_0_135 (.A1(n_0_0_205), .A2(n_0_0_181), .A3(n_0_0_156), .A4(
      n_0_0_131), .ZN(n_0_0_130));
   AOI21_X1 i_0_0_136 (.A(n_0_0_132), .B1(Arr8[15]), .B2(n_0_0_357), .ZN(
      n_0_0_131));
   NAND2_X1 i_0_0_137 (.A1(n_0_0_133), .A2(n_0_0_312), .ZN(n_0_0_132));
   OAI211_X1 i_0_0_138 (.A(n_0_0_135), .B(n_0_0_134), .C1(n_0_0_357), .C2(
      Arr8[15]), .ZN(n_0_0_133));
   NAND2_X1 i_0_0_139 (.A1(n_0_0_356), .A2(Arr8[14]), .ZN(n_0_0_134));
   OAI221_X1 i_0_0_140 (.A(n_0_0_136), .B1(Arr8[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr8[14]), .ZN(n_0_0_135));
   NAND2_X1 i_0_0_141 (.A1(n_0_0_138), .A2(n_0_0_137), .ZN(n_0_0_136));
   AOI22_X1 i_0_0_142 (.A1(n_0_0_355), .A2(Arr8[13]), .B1(n_0_0_354), .B2(
      Arr8[12]), .ZN(n_0_0_137));
   OAI221_X1 i_0_0_143 (.A(n_0_0_139), .B1(Arr8[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr8[12]), .ZN(n_0_0_138));
   NAND2_X1 i_0_0_144 (.A1(n_0_0_141), .A2(n_0_0_140), .ZN(n_0_0_139));
   AOI22_X1 i_0_0_145 (.A1(n_0_0_353), .A2(Arr8[11]), .B1(n_0_0_352), .B2(
      Arr8[10]), .ZN(n_0_0_140));
   OAI221_X1 i_0_0_146 (.A(n_0_0_142), .B1(Arr8[9]), .B2(n_0_0_351), .C1(
      n_0_0_352), .C2(Arr8[10]), .ZN(n_0_0_141));
   NAND2_X1 i_0_0_147 (.A1(n_0_0_144), .A2(n_0_0_143), .ZN(n_0_0_142));
   AOI22_X1 i_0_0_148 (.A1(n_0_0_351), .A2(Arr8[9]), .B1(n_0_0_350), .B2(Arr8[8]), 
      .ZN(n_0_0_143));
   OAI221_X1 i_0_0_149 (.A(n_0_0_145), .B1(Arr8[7]), .B2(n_0_0_349), .C1(
      n_0_0_350), .C2(Arr8[8]), .ZN(n_0_0_144));
   NAND2_X1 i_0_0_150 (.A1(n_0_0_147), .A2(n_0_0_146), .ZN(n_0_0_145));
   AOI22_X1 i_0_0_151 (.A1(n_0_0_349), .A2(Arr8[7]), .B1(n_0_0_348), .B2(Arr8[6]), 
      .ZN(n_0_0_146));
   OAI221_X1 i_0_0_152 (.A(n_0_0_148), .B1(Arr8[5]), .B2(n_0_0_347), .C1(
      n_0_0_348), .C2(Arr8[6]), .ZN(n_0_0_147));
   NAND2_X1 i_0_0_153 (.A1(n_0_0_150), .A2(n_0_0_149), .ZN(n_0_0_148));
   AOI22_X1 i_0_0_154 (.A1(n_0_0_347), .A2(Arr8[5]), .B1(n_0_0_346), .B2(Arr8[4]), 
      .ZN(n_0_0_149));
   OAI21_X1 i_0_0_155 (.A(n_0_0_151), .B1(Arr8[4]), .B2(n_0_0_346), .ZN(
      n_0_0_150));
   OAI21_X1 i_0_0_156 (.A(n_0_0_152), .B1(n_0_0_339), .B2(max[3]), .ZN(n_0_0_151));
   OAI221_X1 i_0_0_157 (.A(n_0_0_153), .B1(Arr8[2]), .B2(n_0_0_344), .C1(
      n_0_0_345), .C2(Arr8[3]), .ZN(n_0_0_152));
   NAND2_X1 i_0_0_158 (.A1(n_0_0_154), .A2(n_0_0_155), .ZN(n_0_0_153));
   AOI22_X1 i_0_0_159 (.A1(n_0_0_344), .A2(Arr8[2]), .B1(n_0_0_343), .B2(Arr8[1]), 
      .ZN(n_0_0_154));
   OAI211_X1 i_0_0_160 (.A(n_0_0_342), .B(Arr8[0]), .C1(n_0_0_343), .C2(Arr8[1]), 
      .ZN(n_0_0_155));
   AOI21_X1 i_0_0_161 (.A(n_0_0_157), .B1(Arr7[15]), .B2(n_0_0_357), .ZN(
      n_0_0_156));
   NAND2_X1 i_0_0_162 (.A1(n_0_0_158), .A2(n_0_0_317), .ZN(n_0_0_157));
   OAI211_X1 i_0_0_163 (.A(n_0_0_160), .B(n_0_0_159), .C1(n_0_0_357), .C2(
      Arr7[15]), .ZN(n_0_0_158));
   NAND2_X1 i_0_0_164 (.A1(n_0_0_356), .A2(Arr7[14]), .ZN(n_0_0_159));
   OAI221_X1 i_0_0_165 (.A(n_0_0_161), .B1(Arr7[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr7[14]), .ZN(n_0_0_160));
   NAND2_X1 i_0_0_166 (.A1(n_0_0_163), .A2(n_0_0_162), .ZN(n_0_0_161));
   AOI22_X1 i_0_0_167 (.A1(n_0_0_355), .A2(Arr7[13]), .B1(n_0_0_354), .B2(
      Arr7[12]), .ZN(n_0_0_162));
   OAI221_X1 i_0_0_168 (.A(n_0_0_164), .B1(Arr7[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr7[12]), .ZN(n_0_0_163));
   NAND2_X1 i_0_0_169 (.A1(n_0_0_166), .A2(n_0_0_165), .ZN(n_0_0_164));
   AOI22_X1 i_0_0_170 (.A1(n_0_0_353), .A2(Arr7[11]), .B1(n_0_0_352), .B2(
      Arr7[10]), .ZN(n_0_0_165));
   OAI221_X1 i_0_0_171 (.A(n_0_0_167), .B1(Arr7[9]), .B2(n_0_0_351), .C1(
      n_0_0_352), .C2(Arr7[10]), .ZN(n_0_0_166));
   NAND2_X1 i_0_0_172 (.A1(n_0_0_169), .A2(n_0_0_168), .ZN(n_0_0_167));
   AOI22_X1 i_0_0_173 (.A1(n_0_0_351), .A2(Arr7[9]), .B1(n_0_0_350), .B2(Arr7[8]), 
      .ZN(n_0_0_168));
   OAI221_X1 i_0_0_174 (.A(n_0_0_170), .B1(Arr7[7]), .B2(n_0_0_349), .C1(
      n_0_0_350), .C2(Arr7[8]), .ZN(n_0_0_169));
   NAND2_X1 i_0_0_175 (.A1(n_0_0_172), .A2(n_0_0_171), .ZN(n_0_0_170));
   AOI22_X1 i_0_0_176 (.A1(n_0_0_349), .A2(Arr7[7]), .B1(n_0_0_348), .B2(Arr7[6]), 
      .ZN(n_0_0_171));
   OAI21_X1 i_0_0_177 (.A(n_0_0_173), .B1(Arr7[6]), .B2(n_0_0_348), .ZN(
      n_0_0_172));
   OAI21_X1 i_0_0_178 (.A(n_0_0_174), .B1(n_0_0_338), .B2(max[5]), .ZN(n_0_0_173));
   OAI221_X1 i_0_0_179 (.A(n_0_0_175), .B1(Arr7[4]), .B2(n_0_0_346), .C1(
      n_0_0_347), .C2(Arr7[5]), .ZN(n_0_0_174));
   NAND2_X1 i_0_0_180 (.A1(n_0_0_177), .A2(n_0_0_176), .ZN(n_0_0_175));
   AOI22_X1 i_0_0_181 (.A1(n_0_0_346), .A2(Arr7[4]), .B1(n_0_0_345), .B2(Arr7[3]), 
      .ZN(n_0_0_176));
   OAI221_X1 i_0_0_182 (.A(n_0_0_178), .B1(Arr7[2]), .B2(n_0_0_344), .C1(
      n_0_0_345), .C2(Arr7[3]), .ZN(n_0_0_177));
   NAND2_X1 i_0_0_183 (.A1(n_0_0_179), .A2(n_0_0_180), .ZN(n_0_0_178));
   AOI22_X1 i_0_0_184 (.A1(n_0_0_344), .A2(Arr7[2]), .B1(n_0_0_343), .B2(Arr7[1]), 
      .ZN(n_0_0_179));
   OAI211_X1 i_0_0_185 (.A(n_0_0_342), .B(Arr7[0]), .C1(n_0_0_343), .C2(Arr7[1]), 
      .ZN(n_0_0_180));
   AOI21_X1 i_0_0_186 (.A(n_0_0_182), .B1(n_0_0_184), .B2(n_0_0_183), .ZN(
      n_0_0_181));
   OAI21_X1 i_0_0_187 (.A(n_0_0_308), .B1(n_0_0_341), .B2(max[15]), .ZN(
      n_0_0_182));
   AOI22_X1 i_0_0_188 (.A1(n_0_0_356), .A2(Arr9[14]), .B1(n_0_0_341), .B2(
      max[15]), .ZN(n_0_0_183));
   OAI221_X1 i_0_0_189 (.A(n_0_0_185), .B1(Arr9[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr9[14]), .ZN(n_0_0_184));
   NAND2_X1 i_0_0_190 (.A1(n_0_0_187), .A2(n_0_0_186), .ZN(n_0_0_185));
   AOI22_X1 i_0_0_191 (.A1(n_0_0_355), .A2(Arr9[13]), .B1(n_0_0_354), .B2(
      Arr9[12]), .ZN(n_0_0_186));
   OAI221_X1 i_0_0_192 (.A(n_0_0_188), .B1(Arr9[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr9[12]), .ZN(n_0_0_187));
   NAND2_X1 i_0_0_193 (.A1(n_0_0_190), .A2(n_0_0_189), .ZN(n_0_0_188));
   AOI22_X1 i_0_0_194 (.A1(n_0_0_353), .A2(Arr9[11]), .B1(n_0_0_352), .B2(
      Arr9[10]), .ZN(n_0_0_189));
   OAI221_X1 i_0_0_195 (.A(n_0_0_191), .B1(Arr9[9]), .B2(n_0_0_351), .C1(
      n_0_0_352), .C2(Arr9[10]), .ZN(n_0_0_190));
   NAND2_X1 i_0_0_196 (.A1(n_0_0_193), .A2(n_0_0_192), .ZN(n_0_0_191));
   AOI22_X1 i_0_0_197 (.A1(n_0_0_351), .A2(Arr9[9]), .B1(n_0_0_350), .B2(Arr9[8]), 
      .ZN(n_0_0_192));
   OAI21_X1 i_0_0_198 (.A(n_0_0_194), .B1(Arr9[8]), .B2(n_0_0_350), .ZN(
      n_0_0_193));
   OAI21_X1 i_0_0_199 (.A(n_0_0_195), .B1(n_0_0_340), .B2(max[7]), .ZN(n_0_0_194));
   OAI221_X1 i_0_0_200 (.A(n_0_0_196), .B1(Arr9[6]), .B2(n_0_0_348), .C1(
      n_0_0_349), .C2(Arr9[7]), .ZN(n_0_0_195));
   NAND2_X1 i_0_0_201 (.A1(n_0_0_198), .A2(n_0_0_197), .ZN(n_0_0_196));
   AOI22_X1 i_0_0_202 (.A1(n_0_0_348), .A2(Arr9[6]), .B1(n_0_0_347), .B2(Arr9[5]), 
      .ZN(n_0_0_197));
   OAI221_X1 i_0_0_203 (.A(n_0_0_199), .B1(Arr9[4]), .B2(n_0_0_346), .C1(
      n_0_0_347), .C2(Arr9[5]), .ZN(n_0_0_198));
   NAND2_X1 i_0_0_204 (.A1(n_0_0_201), .A2(n_0_0_200), .ZN(n_0_0_199));
   AOI22_X1 i_0_0_205 (.A1(n_0_0_346), .A2(Arr9[4]), .B1(n_0_0_345), .B2(Arr9[3]), 
      .ZN(n_0_0_200));
   OAI221_X1 i_0_0_206 (.A(n_0_0_202), .B1(Arr9[2]), .B2(n_0_0_344), .C1(
      n_0_0_345), .C2(Arr9[3]), .ZN(n_0_0_201));
   NAND2_X1 i_0_0_207 (.A1(n_0_0_203), .A2(n_0_0_204), .ZN(n_0_0_202));
   AOI22_X1 i_0_0_208 (.A1(n_0_0_344), .A2(Arr9[2]), .B1(n_0_0_343), .B2(Arr9[1]), 
      .ZN(n_0_0_203));
   OAI211_X1 i_0_0_209 (.A(n_0_0_342), .B(Arr9[0]), .C1(n_0_0_343), .C2(Arr9[1]), 
      .ZN(n_0_0_204));
   AOI21_X1 i_0_0_210 (.A(n_0_0_206), .B1(n_0_0_208), .B2(n_0_0_207), .ZN(
      n_0_0_205));
   OAI21_X1 i_0_0_211 (.A(n_0_0_319), .B1(n_0_0_330), .B2(max[15]), .ZN(
      n_0_0_206));
   AOI22_X1 i_0_0_212 (.A1(n_0_0_356), .A2(Arr2[14]), .B1(n_0_0_330), .B2(
      max[15]), .ZN(n_0_0_207));
   OAI221_X1 i_0_0_213 (.A(n_0_0_209), .B1(Arr2[13]), .B2(n_0_0_355), .C1(
      n_0_0_356), .C2(Arr2[14]), .ZN(n_0_0_208));
   NAND2_X1 i_0_0_214 (.A1(n_0_0_211), .A2(n_0_0_210), .ZN(n_0_0_209));
   AOI22_X1 i_0_0_215 (.A1(n_0_0_355), .A2(Arr2[13]), .B1(n_0_0_354), .B2(
      Arr2[12]), .ZN(n_0_0_210));
   OAI221_X1 i_0_0_216 (.A(n_0_0_212), .B1(Arr2[11]), .B2(n_0_0_353), .C1(
      n_0_0_354), .C2(Arr2[12]), .ZN(n_0_0_211));
   NAND2_X1 i_0_0_217 (.A1(n_0_0_214), .A2(n_0_0_213), .ZN(n_0_0_212));
   AOI22_X1 i_0_0_218 (.A1(n_0_0_353), .A2(Arr2[11]), .B1(n_0_0_352), .B2(
      Arr2[10]), .ZN(n_0_0_213));
   OAI221_X1 i_0_0_219 (.A(n_0_0_215), .B1(Arr2[9]), .B2(n_0_0_351), .C1(
      n_0_0_352), .C2(Arr2[10]), .ZN(n_0_0_214));
   NAND2_X1 i_0_0_220 (.A1(n_0_0_217), .A2(n_0_0_216), .ZN(n_0_0_215));
   AOI22_X1 i_0_0_221 (.A1(n_0_0_351), .A2(Arr2[9]), .B1(n_0_0_350), .B2(Arr2[8]), 
      .ZN(n_0_0_216));
   OAI221_X1 i_0_0_222 (.A(n_0_0_218), .B1(Arr2[7]), .B2(n_0_0_349), .C1(
      n_0_0_350), .C2(Arr2[8]), .ZN(n_0_0_217));
   NAND2_X1 i_0_0_223 (.A1(n_0_0_220), .A2(n_0_0_219), .ZN(n_0_0_218));
   AOI22_X1 i_0_0_224 (.A1(n_0_0_349), .A2(Arr2[7]), .B1(n_0_0_348), .B2(Arr2[6]), 
      .ZN(n_0_0_219));
   OAI221_X1 i_0_0_225 (.A(n_0_0_221), .B1(Arr2[5]), .B2(n_0_0_347), .C1(
      n_0_0_348), .C2(Arr2[6]), .ZN(n_0_0_220));
   NAND2_X1 i_0_0_226 (.A1(n_0_0_223), .A2(n_0_0_222), .ZN(n_0_0_221));
   AOI22_X1 i_0_0_227 (.A1(n_0_0_347), .A2(Arr2[5]), .B1(n_0_0_346), .B2(Arr2[4]), 
      .ZN(n_0_0_222));
   OAI21_X1 i_0_0_228 (.A(n_0_0_224), .B1(Arr2[4]), .B2(n_0_0_346), .ZN(
      n_0_0_223));
   OAI21_X1 i_0_0_229 (.A(n_0_0_225), .B1(n_0_0_329), .B2(max[3]), .ZN(n_0_0_224));
   OAI221_X1 i_0_0_230 (.A(n_0_0_226), .B1(Arr2[2]), .B2(n_0_0_344), .C1(
      n_0_0_345), .C2(Arr2[3]), .ZN(n_0_0_225));
   NAND2_X1 i_0_0_231 (.A1(n_0_0_227), .A2(n_0_0_228), .ZN(n_0_0_226));
   AOI22_X1 i_0_0_232 (.A1(n_0_0_344), .A2(Arr2[2]), .B1(n_0_0_343), .B2(Arr2[1]), 
      .ZN(n_0_0_227));
   OAI211_X1 i_0_0_233 (.A(n_0_0_342), .B(Arr2[0]), .C1(n_0_0_343), .C2(Arr2[1]), 
      .ZN(n_0_0_228));
   NAND3_X1 i_0_0_234 (.A1(n_0_0_233), .A2(n_0_0_232), .A3(n_0_0_229), .ZN(
      n_0_10));
   AOI221_X1 i_0_0_235 (.A(n_0_0_230), .B1(n_0_0_313), .B2(Arr0[0]), .C1(Arr2[0]), 
      .C2(n_0_0_319), .ZN(n_0_0_229));
   INV_X1 i_0_0_236 (.A(n_0_0_231), .ZN(n_0_0_230));
   AOI22_X1 i_0_0_237 (.A1(Arr9[0]), .A2(n_0_0_308), .B1(n_0_0_307), .B2(Arr1[0]), 
      .ZN(n_0_0_231));
   AOI222_X1 i_0_0_238 (.A1(Arr8[0]), .A2(n_0_0_312), .B1(n_0_0_309), .B2(
      Arr6[0]), .C1(Arr4[0]), .C2(n_0_0_314), .ZN(n_0_0_232));
   AOI222_X1 i_0_0_239 (.A1(Arr7[0]), .A2(n_0_0_317), .B1(n_0_0_316), .B2(
      Arr3[0]), .C1(n_0_0_310), .C2(Arr5[0]), .ZN(n_0_0_233));
   NAND3_X1 i_0_0_240 (.A1(n_0_0_236), .A2(n_0_0_235), .A3(n_0_0_234), .ZN(
      n_0_11));
   AOI222_X1 i_0_0_241 (.A1(Arr2[1]), .A2(n_0_0_319), .B1(n_0_0_316), .B2(
      Arr3[1]), .C1(Arr6[1]), .C2(n_0_0_309), .ZN(n_0_0_234));
   AOI222_X1 i_0_0_242 (.A1(Arr7[1]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Arr0[1]), .C1(n_0_0_312), .C2(Arr8[1]), .ZN(n_0_0_235));
   AOI221_X1 i_0_0_243 (.A(n_0_0_237), .B1(n_0_0_307), .B2(Arr1[1]), .C1(Arr9[1]), 
      .C2(n_0_0_308), .ZN(n_0_0_236));
   INV_X1 i_0_0_244 (.A(n_0_0_238), .ZN(n_0_0_237));
   AOI22_X1 i_0_0_245 (.A1(Arr4[1]), .A2(n_0_0_314), .B1(n_0_0_310), .B2(Arr5[1]), 
      .ZN(n_0_0_238));
   NAND3_X1 i_0_0_246 (.A1(n_0_0_241), .A2(n_0_0_240), .A3(n_0_0_239), .ZN(
      n_0_12));
   AOI222_X1 i_0_0_247 (.A1(Arr4[2]), .A2(n_0_0_314), .B1(n_0_0_307), .B2(
      Arr1[2]), .C1(n_0_0_310), .C2(Arr5[2]), .ZN(n_0_0_239));
   AOI222_X1 i_0_0_248 (.A1(Arr2[2]), .A2(n_0_0_319), .B1(n_0_0_309), .B2(
      Arr6[2]), .C1(Arr9[2]), .C2(n_0_0_308), .ZN(n_0_0_240));
   AOI221_X1 i_0_0_249 (.A(n_0_0_242), .B1(n_0_0_316), .B2(Arr3[2]), .C1(Arr8[2]), 
      .C2(n_0_0_312), .ZN(n_0_0_241));
   INV_X1 i_0_0_250 (.A(n_0_0_243), .ZN(n_0_0_242));
   AOI22_X1 i_0_0_251 (.A1(Arr7[2]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(Arr0[2]), 
      .ZN(n_0_0_243));
   NAND3_X1 i_0_0_252 (.A1(n_0_0_248), .A2(n_0_0_247), .A3(n_0_0_244), .ZN(
      n_0_13));
   AOI221_X1 i_0_0_253 (.A(n_0_0_245), .B1(n_0_0_310), .B2(Arr5[3]), .C1(Arr6[3]), 
      .C2(n_0_0_309), .ZN(n_0_0_244));
   INV_X1 i_0_0_254 (.A(n_0_0_246), .ZN(n_0_0_245));
   AOI22_X1 i_0_0_255 (.A1(Arr9[3]), .A2(n_0_0_308), .B1(n_0_0_307), .B2(Arr1[3]), 
      .ZN(n_0_0_246));
   AOI222_X1 i_0_0_256 (.A1(Arr4[3]), .A2(n_0_0_314), .B1(n_0_0_313), .B2(
      Arr0[3]), .C1(n_0_0_312), .C2(Arr8[3]), .ZN(n_0_0_247));
   AOI222_X1 i_0_0_257 (.A1(Arr7[3]), .A2(n_0_0_317), .B1(n_0_0_316), .B2(
      Arr3[3]), .C1(Arr2[3]), .C2(n_0_0_319), .ZN(n_0_0_248));
   NAND3_X1 i_0_0_258 (.A1(n_0_0_251), .A2(n_0_0_250), .A3(n_0_0_249), .ZN(
      n_0_14));
   AOI222_X1 i_0_0_259 (.A1(Arr4[4]), .A2(n_0_0_314), .B1(n_0_0_307), .B2(
      Arr1[4]), .C1(n_0_0_310), .C2(Arr5[4]), .ZN(n_0_0_249));
   AOI222_X1 i_0_0_260 (.A1(Arr2[4]), .A2(n_0_0_319), .B1(n_0_0_309), .B2(
      Arr6[4]), .C1(Arr9[4]), .C2(n_0_0_308), .ZN(n_0_0_250));
   AOI221_X1 i_0_0_261 (.A(n_0_0_252), .B1(n_0_0_316), .B2(Arr3[4]), .C1(Arr8[4]), 
      .C2(n_0_0_312), .ZN(n_0_0_251));
   INV_X1 i_0_0_262 (.A(n_0_0_253), .ZN(n_0_0_252));
   AOI22_X1 i_0_0_263 (.A1(Arr7[4]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(Arr0[4]), 
      .ZN(n_0_0_253));
   NAND3_X1 i_0_0_264 (.A1(n_0_0_256), .A2(n_0_0_255), .A3(n_0_0_254), .ZN(
      n_0_15));
   AOI222_X1 i_0_0_265 (.A1(Arr4[5]), .A2(n_0_0_314), .B1(n_0_0_307), .B2(
      Arr1[5]), .C1(n_0_0_310), .C2(Arr5[5]), .ZN(n_0_0_254));
   AOI222_X1 i_0_0_266 (.A1(Arr2[5]), .A2(n_0_0_319), .B1(n_0_0_309), .B2(
      Arr6[5]), .C1(Arr9[5]), .C2(n_0_0_308), .ZN(n_0_0_255));
   AOI221_X1 i_0_0_267 (.A(n_0_0_257), .B1(n_0_0_316), .B2(Arr3[5]), .C1(Arr8[5]), 
      .C2(n_0_0_312), .ZN(n_0_0_256));
   INV_X1 i_0_0_268 (.A(n_0_0_258), .ZN(n_0_0_257));
   AOI22_X1 i_0_0_269 (.A1(Arr7[5]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(Arr0[5]), 
      .ZN(n_0_0_258));
   NAND3_X1 i_0_0_270 (.A1(n_0_0_261), .A2(n_0_0_260), .A3(n_0_0_259), .ZN(
      n_0_16));
   AOI222_X1 i_0_0_271 (.A1(Arr2[6]), .A2(n_0_0_319), .B1(n_0_0_316), .B2(
      Arr3[6]), .C1(Arr6[6]), .C2(n_0_0_309), .ZN(n_0_0_259));
   AOI222_X1 i_0_0_272 (.A1(Arr7[6]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Arr0[6]), .C1(n_0_0_312), .C2(Arr8[6]), .ZN(n_0_0_260));
   AOI221_X1 i_0_0_273 (.A(n_0_0_262), .B1(n_0_0_307), .B2(Arr1[6]), .C1(Arr9[6]), 
      .C2(n_0_0_308), .ZN(n_0_0_261));
   INV_X1 i_0_0_274 (.A(n_0_0_263), .ZN(n_0_0_262));
   AOI22_X1 i_0_0_275 (.A1(Arr4[6]), .A2(n_0_0_314), .B1(n_0_0_310), .B2(Arr5[6]), 
      .ZN(n_0_0_263));
   NAND3_X1 i_0_0_276 (.A1(n_0_0_266), .A2(n_0_0_265), .A3(n_0_0_264), .ZN(
      n_0_17));
   AOI222_X1 i_0_0_277 (.A1(Arr4[7]), .A2(n_0_0_314), .B1(n_0_0_307), .B2(
      Arr1[7]), .C1(n_0_0_310), .C2(Arr5[7]), .ZN(n_0_0_264));
   AOI222_X1 i_0_0_278 (.A1(Arr2[7]), .A2(n_0_0_319), .B1(n_0_0_309), .B2(
      Arr6[7]), .C1(Arr9[7]), .C2(n_0_0_308), .ZN(n_0_0_265));
   AOI221_X1 i_0_0_279 (.A(n_0_0_267), .B1(n_0_0_316), .B2(Arr3[7]), .C1(Arr8[7]), 
      .C2(n_0_0_312), .ZN(n_0_0_266));
   INV_X1 i_0_0_280 (.A(n_0_0_268), .ZN(n_0_0_267));
   AOI22_X1 i_0_0_281 (.A1(Arr7[7]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(Arr0[7]), 
      .ZN(n_0_0_268));
   NAND3_X1 i_0_0_282 (.A1(n_0_0_273), .A2(n_0_0_272), .A3(n_0_0_269), .ZN(
      n_0_18));
   AOI221_X1 i_0_0_283 (.A(n_0_0_270), .B1(n_0_0_313), .B2(Arr0[8]), .C1(Arr2[8]), 
      .C2(n_0_0_319), .ZN(n_0_0_269));
   INV_X1 i_0_0_284 (.A(n_0_0_271), .ZN(n_0_0_270));
   AOI22_X1 i_0_0_285 (.A1(Arr9[8]), .A2(n_0_0_308), .B1(n_0_0_307), .B2(Arr1[8]), 
      .ZN(n_0_0_271));
   AOI222_X1 i_0_0_286 (.A1(Arr8[8]), .A2(n_0_0_312), .B1(n_0_0_309), .B2(
      Arr6[8]), .C1(Arr4[8]), .C2(n_0_0_314), .ZN(n_0_0_272));
   AOI222_X1 i_0_0_287 (.A1(Arr7[8]), .A2(n_0_0_317), .B1(n_0_0_316), .B2(
      Arr3[8]), .C1(n_0_0_310), .C2(Arr5[8]), .ZN(n_0_0_273));
   NAND3_X1 i_0_0_288 (.A1(n_0_0_276), .A2(n_0_0_275), .A3(n_0_0_274), .ZN(
      n_0_19));
   AOI222_X1 i_0_0_289 (.A1(Arr2[9]), .A2(n_0_0_319), .B1(n_0_0_316), .B2(
      Arr3[9]), .C1(Arr6[9]), .C2(n_0_0_309), .ZN(n_0_0_274));
   AOI222_X1 i_0_0_290 (.A1(Arr7[9]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Arr0[9]), .C1(n_0_0_312), .C2(Arr8[9]), .ZN(n_0_0_275));
   AOI221_X1 i_0_0_291 (.A(n_0_0_277), .B1(n_0_0_307), .B2(Arr1[9]), .C1(Arr9[9]), 
      .C2(n_0_0_308), .ZN(n_0_0_276));
   INV_X1 i_0_0_292 (.A(n_0_0_278), .ZN(n_0_0_277));
   AOI22_X1 i_0_0_293 (.A1(Arr4[9]), .A2(n_0_0_314), .B1(n_0_0_310), .B2(Arr5[9]), 
      .ZN(n_0_0_278));
   NAND3_X1 i_0_0_294 (.A1(n_0_0_283), .A2(n_0_0_282), .A3(n_0_0_279), .ZN(
      n_0_20));
   AOI221_X1 i_0_0_295 (.A(n_0_0_280), .B1(n_0_0_313), .B2(Arr0[10]), .C1(
      Arr2[10]), .C2(n_0_0_319), .ZN(n_0_0_279));
   INV_X1 i_0_0_296 (.A(n_0_0_281), .ZN(n_0_0_280));
   AOI22_X1 i_0_0_297 (.A1(Arr9[10]), .A2(n_0_0_308), .B1(n_0_0_307), .B2(
      Arr1[10]), .ZN(n_0_0_281));
   AOI222_X1 i_0_0_298 (.A1(Arr8[10]), .A2(n_0_0_312), .B1(n_0_0_309), .B2(
      Arr6[10]), .C1(Arr4[10]), .C2(n_0_0_314), .ZN(n_0_0_282));
   AOI222_X1 i_0_0_299 (.A1(Arr7[10]), .A2(n_0_0_317), .B1(n_0_0_316), .B2(
      Arr3[10]), .C1(n_0_0_310), .C2(Arr5[10]), .ZN(n_0_0_283));
   NAND3_X1 i_0_0_300 (.A1(n_0_0_286), .A2(n_0_0_285), .A3(n_0_0_284), .ZN(
      n_0_21));
   AOI222_X1 i_0_0_301 (.A1(Arr2[11]), .A2(n_0_0_319), .B1(n_0_0_316), .B2(
      Arr3[11]), .C1(Arr6[11]), .C2(n_0_0_309), .ZN(n_0_0_284));
   AOI222_X1 i_0_0_302 (.A1(Arr7[11]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Arr0[11]), .C1(n_0_0_312), .C2(Arr8[11]), .ZN(n_0_0_285));
   AOI221_X1 i_0_0_303 (.A(n_0_0_287), .B1(n_0_0_307), .B2(Arr1[11]), .C1(
      Arr9[11]), .C2(n_0_0_308), .ZN(n_0_0_286));
   INV_X1 i_0_0_304 (.A(n_0_0_288), .ZN(n_0_0_287));
   AOI22_X1 i_0_0_305 (.A1(Arr4[11]), .A2(n_0_0_314), .B1(n_0_0_310), .B2(
      Arr5[11]), .ZN(n_0_0_288));
   NAND3_X1 i_0_0_306 (.A1(n_0_0_291), .A2(n_0_0_290), .A3(n_0_0_289), .ZN(
      n_0_22));
   AOI222_X1 i_0_0_307 (.A1(Arr4[12]), .A2(n_0_0_314), .B1(n_0_0_307), .B2(
      Arr1[12]), .C1(n_0_0_310), .C2(Arr5[12]), .ZN(n_0_0_289));
   AOI222_X1 i_0_0_308 (.A1(Arr2[12]), .A2(n_0_0_319), .B1(n_0_0_309), .B2(
      Arr6[12]), .C1(Arr9[12]), .C2(n_0_0_308), .ZN(n_0_0_290));
   AOI221_X1 i_0_0_309 (.A(n_0_0_292), .B1(n_0_0_316), .B2(Arr3[12]), .C1(
      Arr8[12]), .C2(n_0_0_312), .ZN(n_0_0_291));
   INV_X1 i_0_0_310 (.A(n_0_0_293), .ZN(n_0_0_292));
   AOI22_X1 i_0_0_311 (.A1(Arr7[12]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Arr0[12]), .ZN(n_0_0_293));
   NAND3_X1 i_0_0_312 (.A1(n_0_0_296), .A2(n_0_0_295), .A3(n_0_0_294), .ZN(
      n_0_23));
   AOI222_X1 i_0_0_313 (.A1(Arr4[13]), .A2(n_0_0_314), .B1(n_0_0_307), .B2(
      Arr1[13]), .C1(n_0_0_310), .C2(Arr5[13]), .ZN(n_0_0_294));
   AOI222_X1 i_0_0_314 (.A1(Arr2[13]), .A2(n_0_0_319), .B1(n_0_0_309), .B2(
      Arr6[13]), .C1(Arr9[13]), .C2(n_0_0_308), .ZN(n_0_0_295));
   AOI221_X1 i_0_0_315 (.A(n_0_0_297), .B1(n_0_0_316), .B2(Arr3[13]), .C1(
      Arr8[13]), .C2(n_0_0_312), .ZN(n_0_0_296));
   INV_X1 i_0_0_316 (.A(n_0_0_298), .ZN(n_0_0_297));
   AOI22_X1 i_0_0_317 (.A1(Arr7[13]), .A2(n_0_0_317), .B1(n_0_0_313), .B2(
      Arr0[13]), .ZN(n_0_0_298));
   NAND3_X1 i_0_0_318 (.A1(n_0_0_303), .A2(n_0_0_302), .A3(n_0_0_299), .ZN(
      n_0_24));
   AOI221_X1 i_0_0_319 (.A(n_0_0_300), .B1(n_0_0_310), .B2(Arr5[14]), .C1(
      Arr6[14]), .C2(n_0_0_309), .ZN(n_0_0_299));
   INV_X1 i_0_0_320 (.A(n_0_0_301), .ZN(n_0_0_300));
   AOI22_X1 i_0_0_321 (.A1(Arr9[14]), .A2(n_0_0_308), .B1(n_0_0_307), .B2(
      Arr1[14]), .ZN(n_0_0_301));
   AOI222_X1 i_0_0_322 (.A1(Arr4[14]), .A2(n_0_0_314), .B1(n_0_0_313), .B2(
      Arr0[14]), .C1(n_0_0_312), .C2(Arr8[14]), .ZN(n_0_0_302));
   AOI222_X1 i_0_0_323 (.A1(Arr7[14]), .A2(n_0_0_317), .B1(n_0_0_316), .B2(
      Arr3[14]), .C1(Arr2[14]), .C2(n_0_0_319), .ZN(n_0_0_303));
   NAND3_X1 i_0_0_324 (.A1(n_0_0_315), .A2(n_0_0_311), .A3(n_0_0_304), .ZN(
      n_0_25));
   AOI221_X1 i_0_0_325 (.A(n_0_0_305), .B1(n_0_0_310), .B2(Arr5[15]), .C1(
      Arr6[15]), .C2(n_0_0_309), .ZN(n_0_0_304));
   INV_X1 i_0_0_326 (.A(n_0_0_306), .ZN(n_0_0_305));
   AOI22_X1 i_0_0_327 (.A1(Arr9[15]), .A2(n_0_0_308), .B1(n_0_0_307), .B2(
      Arr1[15]), .ZN(n_0_0_306));
   NOR3_X1 i_0_0_328 (.A1(n_0_6), .A2(i[3]), .A3(n_0_0_325), .ZN(n_0_0_307));
   NOR3_X1 i_0_0_329 (.A1(n_0_0_327), .A2(n_0_0_325), .A3(n_0_0_322), .ZN(
      n_0_0_308));
   AND3_X1 i_0_0_330 (.A1(i[2]), .A2(maxIndex[1]), .A3(n_0_0_327), .ZN(n_0_0_309));
   NOR3_X1 i_0_0_331 (.A1(n_0_0_318), .A2(i[1]), .A3(n_0_0_327), .ZN(n_0_0_310));
   NAND2_X1 i_0_0_332 (.A1(i[0]), .A2(n_0_0_323), .ZN(n_0_6));
   AOI222_X1 i_0_0_333 (.A1(Arr4[15]), .A2(n_0_0_314), .B1(n_0_0_313), .B2(
      Arr0[15]), .C1(n_0_0_312), .C2(Arr8[15]), .ZN(n_0_0_311));
   NOR2_X1 i_0_0_334 (.A1(n_0_0_324), .A2(n_0_0_322), .ZN(n_0_0_312));
   AOI21_X1 i_0_0_335 (.A(maxIndex[3]), .B1(n_0_0_324), .B2(n_0_0_321), .ZN(
      n_0_0_313));
   NOR2_X1 i_0_0_336 (.A1(n_0_0_325), .A2(n_0_0_322), .ZN(maxIndex[3]));
   NOR3_X1 i_0_0_337 (.A1(n_0_0_318), .A2(i[0]), .A3(i[1]), .ZN(n_0_0_314));
   AOI222_X1 i_0_0_338 (.A1(Arr7[15]), .A2(n_0_0_317), .B1(n_0_0_316), .B2(
      Arr3[15]), .C1(Arr2[15]), .C2(n_0_0_319), .ZN(n_0_0_315));
   NOR3_X1 i_0_0_339 (.A1(n_0_0_320), .A2(i[2]), .A3(n_0_0_327), .ZN(n_0_0_316));
   AND3_X1 i_0_0_340 (.A1(i[2]), .A2(i[0]), .A3(maxIndex[1]), .ZN(n_0_0_317));
   INV_X1 i_0_0_341 (.A(n_0_0_318), .ZN(maxIndex[2]));
   NAND2_X1 i_0_0_342 (.A1(i[2]), .A2(n_0_0_321), .ZN(n_0_0_318));
   NOR3_X1 i_0_0_343 (.A1(n_0_0_320), .A2(i[0]), .A3(i[2]), .ZN(n_0_0_319));
   INV_X1 i_0_0_344 (.A(n_0_0_320), .ZN(maxIndex[1]));
   NAND2_X1 i_0_0_345 (.A1(i[1]), .A2(n_0_0_321), .ZN(n_0_0_320));
   NOR3_X1 i_0_0_346 (.A1(n_0_0_326), .A2(done), .A3(i[3]), .ZN(n_0_0_321));
   AND3_X1 i_0_0_347 (.A1(n_0_0_324), .A2(n_0_0_323), .A3(i[3]), .ZN(n_0_26));
   NAND2_X1 i_0_0_348 (.A1(i[3]), .A2(n_0_0_323), .ZN(n_0_0_322));
   NOR2_X1 i_0_0_349 (.A1(n_0_0_326), .A2(done), .ZN(n_0_0_323));
   OR2_X1 i_0_0_350 (.A1(n_0_0_325), .A2(i[0]), .ZN(n_0_0_324));
   OR2_X1 i_0_0_351 (.A1(i[2]), .A2(i[1]), .ZN(n_0_0_325));
   INV_X1 i_0_0_352 (.A(enable), .ZN(n_0_0_326));
   INV_X1 i_0_0_353 (.A(i[0]), .ZN(n_0_0_327));
   INV_X1 i_0_0_354 (.A(Arr1[9]), .ZN(n_0_0_328));
   INV_X1 i_0_0_355 (.A(Arr2[3]), .ZN(n_0_0_329));
   INV_X1 i_0_0_356 (.A(Arr2[15]), .ZN(n_0_0_330));
   INV_X1 i_0_0_357 (.A(Arr3[3]), .ZN(n_0_0_331));
   INV_X1 i_0_0_358 (.A(Arr3[15]), .ZN(n_0_0_332));
   INV_X1 i_0_0_359 (.A(Arr4[3]), .ZN(n_0_0_333));
   INV_X1 i_0_0_360 (.A(Arr4[15]), .ZN(n_0_0_334));
   INV_X1 i_0_0_361 (.A(Arr5[7]), .ZN(n_0_0_335));
   INV_X1 i_0_0_362 (.A(Arr5[15]), .ZN(n_0_0_336));
   INV_X1 i_0_0_363 (.A(Arr6[3]), .ZN(n_0_0_337));
   INV_X1 i_0_0_364 (.A(Arr7[5]), .ZN(n_0_0_338));
   INV_X1 i_0_0_365 (.A(Arr8[3]), .ZN(n_0_0_339));
   INV_X1 i_0_0_366 (.A(Arr9[7]), .ZN(n_0_0_340));
   INV_X1 i_0_0_367 (.A(Arr9[15]), .ZN(n_0_0_341));
   INV_X1 i_0_0_368 (.A(max[0]), .ZN(n_0_0_342));
   INV_X1 i_0_0_369 (.A(max[1]), .ZN(n_0_0_343));
   INV_X1 i_0_0_370 (.A(max[2]), .ZN(n_0_0_344));
   INV_X1 i_0_0_371 (.A(max[3]), .ZN(n_0_0_345));
   INV_X1 i_0_0_372 (.A(max[4]), .ZN(n_0_0_346));
   INV_X1 i_0_0_373 (.A(max[5]), .ZN(n_0_0_347));
   INV_X1 i_0_0_374 (.A(max[6]), .ZN(n_0_0_348));
   INV_X1 i_0_0_375 (.A(max[7]), .ZN(n_0_0_349));
   INV_X1 i_0_0_376 (.A(max[8]), .ZN(n_0_0_350));
   INV_X1 i_0_0_377 (.A(max[9]), .ZN(n_0_0_351));
   INV_X1 i_0_0_378 (.A(max[10]), .ZN(n_0_0_352));
   INV_X1 i_0_0_379 (.A(max[11]), .ZN(n_0_0_353));
   INV_X1 i_0_0_380 (.A(max[12]), .ZN(n_0_0_354));
   INV_X1 i_0_0_381 (.A(max[13]), .ZN(n_0_0_355));
   INV_X1 i_0_0_382 (.A(max[14]), .ZN(n_0_0_356));
   INV_X1 i_0_0_383 (.A(max[15]), .ZN(n_0_0_357));
endmodule
